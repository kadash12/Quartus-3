library ieee;
use ieee.std_logic_1164.all;

entity not_DFF_Traf_Cont is port(
	EV_L,CW: in std_logic;
	Q3,Q2,Q1,Q0: in std_logic;
	D3,J2,K2,J1,K1,T0: out std_logic;
	G,Y,R: out std_logic
);
end not_DFF_Traf_Cont;

architecture logic of not_DFF_Traf_Cont is 
signal EV: std_logic;
begin 
	-- Define inputs
	EV <= not EV_L;
	
	--D3 = (/Q3Q2Q1Q0) + (Q3/Q2/Q1/Q0) + (Q3/Q2/Q1Q0EV)
	D3 <= ((NOT Q3) AND Q2 AND Q1 AND Q0)
	OR (Q3 AND (NOT Q2) AND (NOT Q1) AND (NOT Q0))
	OR (Q3 AND (NOT Q2) AND (NOT Q1) AND Q0 AND EV);
	
	--J2 = (/Q3/Q2/Q1/Q0EV) + (/Q3/Q2/Q1Q0EV) + (/Q3/Q2Q1/Q0EV) + (/Q3/Q2Q1Q0/EV) +
	--		 (/Q3/Q2Q1Q0EV)
	J2 <= ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND (NOT Q0) AND EV)
	OR ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND Q0 AND EV)
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND (NOT Q0) AND EV)
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND Q0 AND EV) 
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND Q0 AND (NOT EV) AND CW);
	
	--K2 = (/Q3Q2/Q1/Q0) + (/Q3Q2Q1Q0)
	K2 <= ((NOT Q3) AND Q2 AND (NOT Q1) AND (NOT Q0) AND (NOT CW))
	OR ((NOT Q3) AND Q2 AND Q1 AND Q0);
	
	--J1 = (/Q3/Q2/Q1/Q0EV) + (/Q3/Q2/Q1Q0/EV) + (/Q3/Q2/Q1Q0EV) + (/Q3Q2/Q1Q0) 
	J1 <= ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND (NOT Q0) AND EV)
	OR ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND Q0 AND (NOT EV))
	OR ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND Q0 AND EV)
	OR ((NOT Q3) AND Q2 AND (NOT Q1) AND Q0);
	
	--K1 = (/Q3/Q2Q1Q0/EV) + (/Q3Q2Q1Q0)
	K1 <= ((NOT Q3) AND (NOT Q2) AND Q1 AND Q0 AND (NOT EV) AND (NOT CW))
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND Q0 AND (NOT EV) AND CW)
	OR ((NOT Q3) AND Q2 AND Q1 AND Q0);
	
	--T = (Q3+Q2+Q1+Q0+/EV) (Q3+Q2+/Q1+Q0+/EV) (Q3+/Q2+Q1+Q0+CW) (/Q3+Q2+Q1+/Q0+/EV)
	T0 <= (Q3 OR Q2 OR Q1 OR Q0 OR (NOT EV)) 
	AND (Q3 OR Q2 OR (NOT Q1) OR Q0 OR (NOT EV)) 
	AND (Q3 OR (NOT Q2) OR Q1 OR Q0 OR CW)
	AND ((NOT Q3) OR Q2 OR Q1 OR (NOT Q0) OR (NOT EV))
	AND (Q3 OR Q2 OR (NOT Q1) OR (NOT Q0) OR EV OR (NOT CW));
	
	--G = (/Q3/Q2/Q1/Q0/EV) + (/Q3/Q2/Q1Q0/EV) + (/Q3/Q2Q1/Q0/EV) + (/Q3/Q2Q1Q0/EV) +
	--		(/Q3Q2/Q1/Q0/CW) + (/Q3Q2/Q1/Q0CW)
	G <= ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND (NOT Q0) AND (NOT EV))
	OR ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND Q0 AND (NOT EV))
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND (NOT Q0) AND (NOT EV))
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND Q0 AND (NOT EV) AND (NOT CW)) 
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND Q0 AND (NOT EV) AND CW)
	OR ((NOT Q3) AND Q2 AND (NOT Q1) AND (NOT Q0) AND (NOT CW))
	OR ((NOT Q3) AND Q2 AND (NOT Q1) AND (NOT Q0) AND CW);

	--Y = (/Q3/Q2/Q1/Q0EV) + (/Q3/Q2/Q1Q0EV) + (/Q3/Q2Q1/Q0EV) + (/Q3/Q2Q1Q0EV) + 
	--	   (/Q3Q2/Q1Q0) + (/Q3Q2Q1/Q0)
	Y <= ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND (NOT Q0) AND EV)
	OR ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND Q0 AND EV)
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND (NOT Q0) AND EV)
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND Q0 AND EV)
	OR ((NOT Q3) AND Q2 AND (NOT Q1) AND Q0)
	OR ((NOT Q3) AND Q2 AND Q1 AND (NOT Q0));
	
	--R = (/Q3Q2Q1Q0) + (Q3/Q2/Q1/Q0) + (Q3/Q2/Q1Q0/EV) + (Q3/Q2/Q1Q0/EV)
	R <= ((NOT Q3) AND Q2 AND Q1 AND Q0)
	OR (Q3 AND (NOT Q2) AND (NOT Q1) AND (NOT Q0))
	OR (Q3 AND (NOT Q2) AND (NOT Q1) AND Q0 AND (NOT EV))
	OR (Q3 AND (NOT Q2) AND (NOT Q1) AND Q0 AND EV);
	
	end logic;