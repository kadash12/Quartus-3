library ieee;
use ieee.std_logic_1164.all;

entity DFF_Traf_Cont is port(
	EV_L,CW: in std_logic;
	Q3,Q2,Q1,Q0: in std_logic;
	D3,D2,D1,D0: out std_logic;
	G,Y,R: out std_logic
);
end DFF_Traf_Cont;

architecture logic of DFF_Traf_Cont is 
signal EV: std_logic;
begin 
	-- Define inputs
	EV <= not EV_L;
	
	--D3 = (/Q3Q2Q1Q0) + (Q3/Q2/Q1/Q0) + (Q3/Q2/Q1Q0EV)
	D3 <= ((NOT Q3) AND Q2 AND Q1 AND Q0)
	OR (Q3 AND (NOT Q2) AND (NOT Q1) AND (NOT Q0))
	OR (Q3 AND (NOT Q2) AND (NOT Q1) AND Q0 AND EV);
	
	--D2 = (/Q3/Q2/Q1/Q0EV) + (/Q3/Q2/Q1Q0EV) + (/Q3/Q2Q1/Q0EV) + (/Q3/Q2Q1Q0/EV) +
	--		 (/Q3/Q2Q1Q0EV) + (/Q3Q2/Q1/Q0CW) + (/Q3Q2/Q1Q0) + (/Q3Q2Q1/Q0)
	D2 <= ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND (NOT Q0) AND EV)
	OR ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND Q0 AND EV)
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND (NOT Q0) AND EV)
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND Q0 AND EV)
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND Q0 AND (NOT EV) AND CW) 
	OR ((NOT Q3) AND Q2 AND (NOT Q1) AND Q0)
	OR ((NOT Q3) AND Q2 AND Q1 AND (NOT Q0));
	
	--D1 = (/Q3/Q2/Q1/Q0EV) + (/Q3/Q2/Q1Q0/EV) + (/Q3/Q2/Q1Q0EV) + (/Q3/Q2Q1/Q0/EV) +
	--		 (/Q3/Q2Q1/Q0EV) + (/Q3/Q2Q1Q0EV) + (/Q3Q2/Q1Q0) + (/Q3Q2Q1/Q0)
	D1 <= ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND (NOT Q0) AND EV)
	OR ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND Q0 AND (NOT EV))
	OR ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND Q0 AND EV)
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND (NOT Q0) AND (NOT EV))
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND (NOT Q0) AND EV)
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND Q0 AND EV)
	OR ((NOT Q3) AND Q2 AND (NOT Q1) AND Q0)
	OR ((NOT Q3) AND Q2 AND Q1 AND (NOT Q0));
	
	--D0 = (/Q3/Q2/Q1/Q0/EV) + (/Q3/Q2Q1/Q0/EV) + (/Q3Q2/Q1/Q0CW) + (/Q3Q2Q1/Q0) + 
	--		 (Q3/Q2/Q1/Q0) + (Q3/Q2/Q1Q0EV)
	D0 <= ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND (NOT Q0) AND (NOT EV))
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND (NOT Q0) AND (NOT EV))
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND Q0 AND (NOT EV) AND CW)
	OR ((NOT Q3) AND Q2 AND Q1 AND (NOT Q0))
	OR (Q3 AND (NOT Q2) AND (NOT Q1) AND (NOT Q0))
	OR (Q3 AND (NOT Q2) AND (NOT Q1) AND Q0 AND EV);
	
	--G = (/Q3/Q2/Q1/Q0/EV) + (/Q3/Q2/Q1Q0/EV) + (/Q3/Q2Q1/Q0/EV) + (/Q3/Q2Q1Q0/EV) +
	--		(/Q3Q2/Q1/Q0/CW) + (/Q3Q2/Q1/Q0CW)
	G <= ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND (NOT Q0) AND (NOT EV))
	OR ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND Q0 AND (NOT EV))
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND (NOT Q0) AND (NOT EV))
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND Q0 AND (NOT EV) AND (NOT CW)) 
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND Q0 AND (NOT EV) AND CW);			

	--Y = (/Q3/Q2/Q1/Q0EV) + (/Q3/Q2/Q1Q0EV) + (/Q3/Q2Q1/Q0EV) + (/Q3/Q2Q1Q0EV) + 
	--	   (/Q3Q2/Q1Q0) + (/Q3Q2Q1/Q0)
	Y <= ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND (NOT Q0) AND EV)
	OR ((NOT Q3) AND (NOT Q2) AND (NOT Q1) AND Q0 AND EV)
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND (NOT Q0) AND EV)
	OR ((NOT Q3) AND (NOT Q2) AND Q1 AND Q0 AND EV)
	OR ((NOT Q3) AND Q2 AND (NOT Q1) AND Q0)
	OR ((NOT Q3) AND Q2 AND Q1 AND (NOT Q0));
	
	--R = (/Q3Q2Q1Q0) + (Q3/Q2/Q1/Q0) + (Q3/Q2/Q1Q0/EV) + (Q3/Q2/Q1Q0/EV)
	R <= ((NOT Q3) AND Q2 AND Q1 AND Q0)
	OR (Q3 AND (NOT Q2) AND (NOT Q1) AND (NOT Q0))
	OR (Q3 AND (NOT Q2) AND (NOT Q1) AND Q0 AND (NOT EV))
	OR (Q3 AND (NOT Q2) AND (NOT Q1) AND Q0 AND EV);
	
	end logic;